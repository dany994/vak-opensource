module top();
    reg [64-1:0] a;
    reg [64-1:0] b;
    reg [64-1:0] c;
    always @(*) b[0] <= ~(a[18] ^ a[27]);
    always @(*) b[1] <= (a[10] | a[9]);
    always @(*) b[2] <= a[42] ^ a[55];
    always @(*) b[3] <= (a[13] | a[53]);
    always @(*) b[4] <= ~(a[0] ^ a[14]);
    always @(*) b[5] <= (a[13] | a[57]);
    always @(*) b[6] <= ~(a[63] ^ a[16]);
    always @(*) b[7] <= ~(a[41] ^ a[26]);
    always @(*) b[8] <= a[31] ^ a[62];
    always @(*) b[9] <= ~(a[18] ^ a[54]);
    always @(*) b[10] <= a[57] & a[5];
    always @(*) b[11] <= ~(a[5] ^ a[50]);
    always @(*) b[12] <= ~(a[28] ^ a[47]);
    always @(*) b[13] <= ~(a[55] | a[6]);
    always @(*) b[14] <= ~(a[24] ^ a[48]);
    always @(*) b[15] <= ~(a[45] ^ a[28]);
    always @(*) b[16] <= ~(a[36] | a[26]);
    always @(*) b[17] <= ~(a[39] & a[55]);
    always @(*) b[18] <= ~(a[26] & a[57]);
    always @(*) b[19] <= a[39] ^ a[32];
    always @(*) b[20] <= ~(a[13] & a[55]);
    always @(*) b[21] <= (a[51] | a[46]);
    always @(*) b[22] <= a[18] ^ a[51];
    always @(*) b[23] <= a[17] ^ a[43];
    always @(*) b[24] <= (a[16] | a[2]);
    always @(*) b[25] <= ~(a[30] | a[32]);
    always @(*) b[26] <= a[44] & a[62];
    always @(*) b[27] <= ~(a[52] ^ a[25]);
    always @(*) b[28] <= ~(a[36] | a[61]);
    always @(*) b[29] <= ~(a[21] | a[48]);
    always @(*) b[30] <= ~(a[47] & a[56]);
    always @(*) b[31] <= ~(a[56] & a[17]);
    always @(*) b[32] <= ~(a[18] ^ a[4]);
    always @(*) b[33] <= ~(a[56] & a[52]);
    always @(*) b[34] <= ~(a[48] ^ a[28]);
    always @(*) b[35] <= a[40] & a[49];
    always @(*) b[36] <= (a[40] | a[5]);
    always @(*) b[37] <= ~(a[7] & a[11]);
    always @(*) b[38] <= a[33] ^ a[28];
    always @(*) b[39] <= a[0] & a[9];
    always @(*) b[40] <= (a[30] | a[24]);
    always @(*) b[41] <= a[38] & a[5];
    always @(*) b[42] <= (a[10] | a[41]);
    always @(*) b[43] <= a[24] & a[39];
    always @(*) b[44] <= a[41] ^ a[54];
    always @(*) b[45] <= ~(a[29] & a[32]);
    always @(*) b[46] <= a[18] & a[54];
    always @(*) b[47] <= ~(a[45] ^ a[55]);
    always @(*) b[48] <= ~(a[15] ^ a[16]);
    always @(*) b[49] <= ~(a[13] & a[55]);
    always @(*) b[50] <= ~(a[28] & a[6]);
    always @(*) b[51] <= ~(a[5] & a[37]);
    always @(*) b[52] <= a[50] & a[42];
    always @(*) b[53] <= ~(a[57] ^ a[5]);
    always @(*) b[54] <= ~(a[35] | a[10]);
    always @(*) b[55] <= a[49] ^ a[38];
    always @(*) b[56] <= ~(a[46] | a[48]);
    always @(*) b[57] <= ~(a[56] | a[33]);
    always @(*) b[58] <= ~(a[55] & a[55]);
    always @(*) b[59] <= a[40] & a[22];
    always @(*) b[60] <= ~(a[14] ^ a[61]);
    always @(*) b[61] <= ~(a[28] ^ a[53]);
    always @(*) b[62] <= (a[49] | a[23]);
    always @(*) b[63] <= ~(a[4] ^ a[11]);
    always @(*) c[0] <= ~(b[20] & b[3]);
    always @(*) c[1] <= ~(b[58] & b[63]);
    always @(*) c[2] <= (b[23] | b[22]);
    always @(*) c[3] <= ~(b[50] | b[25]);
    always @(*) c[4] <= b[39] ^ b[3];
    always @(*) c[5] <= ~(b[57] & b[22]);
    always @(*) c[6] <= b[44] ^ b[9];
    always @(*) c[7] <= ~(b[49] | b[61]);
    always @(*) c[8] <= ~(b[50] | b[9]);
    always @(*) c[9] <= b[10] ^ b[49];
    always @(*) c[10] <= b[63] & b[20];
    always @(*) c[11] <= (b[22] | b[60]);
    always @(*) c[12] <= b[37] ^ b[9];
    always @(*) c[13] <= ~(b[43] ^ b[54]);
    always @(*) c[14] <= ~(b[62] ^ b[43]);
    always @(*) c[15] <= ~(b[63] & b[47]);
    always @(*) c[16] <= b[57] ^ b[44];
    always @(*) c[17] <= ~(b[32] & b[11]);
    always @(*) c[18] <= b[57] ^ b[53];
    always @(*) c[19] <= b[24] ^ b[51];
    always @(*) c[20] <= (b[53] | b[48]);
    always @(*) c[21] <= ~(b[12] ^ b[27]);
    always @(*) c[22] <= b[32] ^ b[4];
    always @(*) c[23] <= ~(b[37] ^ b[2]);
    always @(*) c[24] <= (b[34] | b[4]);
    always @(*) c[25] <= (b[9] | b[24]);
    always @(*) c[26] <= (b[60] | b[13]);
    always @(*) c[27] <= ~(b[22] & b[39]);
    always @(*) c[28] <= ~(b[60] & b[39]);
    always @(*) c[29] <= b[32] ^ b[14];
    always @(*) c[30] <= ~(b[57] | b[49]);
    always @(*) c[31] <= b[61] & b[44];
    always @(*) c[32] <= b[19] ^ b[20];
    always @(*) c[33] <= ~(b[45] ^ b[24]);
    always @(*) c[34] <= ~(b[31] | b[35]);
    always @(*) c[35] <= b[23] ^ b[63];
    always @(*) c[36] <= (b[5] | b[48]);
    always @(*) c[37] <= b[20] ^ b[26];
    always @(*) c[38] <= b[30] ^ b[21];
    always @(*) c[39] <= b[62] & b[54];
    always @(*) c[40] <= b[13] & b[36];
    always @(*) c[41] <= ~(b[37] & b[22]);
    always @(*) c[42] <= ~(b[26] | b[25]);
    always @(*) c[43] <= b[8] & b[18];
    always @(*) c[44] <= ~(b[47] | b[61]);
    always @(*) c[45] <= ~(b[40] | b[15]);
    always @(*) c[46] <= ~(b[11] & b[39]);
    always @(*) c[47] <= ~(b[17] ^ b[61]);
    always @(*) c[48] <= ~(b[15] | b[26]);
    always @(*) c[49] <= ~(b[45] & b[48]);
    always @(*) c[50] <= b[15] & b[44];
    always @(*) c[51] <= ~(b[38] & b[44]);
    always @(*) c[52] <= ~(b[54] | b[13]);
    always @(*) c[53] <= b[37] ^ b[28];
    always @(*) c[54] <= b[61] & b[33];
    always @(*) c[55] <= ~(b[39] ^ b[17]);
    always @(*) c[56] <= (b[20] | b[37]);
    always @(*) c[57] <= ~(b[47] | b[3]);
    always @(*) c[58] <= ~(b[11] ^ b[25]);
    always @(*) c[59] <= b[30] ^ b[50];
    always @(*) c[60] <= ~(b[55] & b[47]);
    always @(*) c[61] <= ~(b[34] & b[30]);
    always @(*) c[62] <= b[56] ^ b[42];
    always @(*) c[63] <= ~(b[20] | b[0]);

    integer i;
    initial begin
        a = 0;
        b = 0;
        c = 0;
        for (i=0; i<400; i=i+1) begin
            a[12] <= ~a[12];
            a[2] <= ~a[2];
            a[3] <= ~a[3];
            #1;
            a[32] <= ~a[32];
            a[56] <= ~a[56];
            a[57] <= ~a[57];
            #1;
            a[28] <= ~a[28];
            a[14] <= ~a[14];
            a[51] <= ~a[51];
            #1;
            a[57] <= ~a[57];
            a[34] <= ~a[34];
            #1;
            a[59] <= ~a[59];
            a[26] <= ~a[26];
            a[48] <= ~a[48];
            a[34] <= ~a[34];
            #1;
            a[19] <= ~a[19];
            a[48] <= ~a[48];
            a[2] <= ~a[2];
            a[35] <= ~a[35];
            a[9] <= ~a[9];
            a[9] <= ~a[9];
            a[28] <= ~a[28];
            a[12] <= ~a[12];
            a[9] <= ~a[9];
            a[37] <= ~a[37];
            a[31] <= ~a[31];
            a[17] <= ~a[17];
            a[8] <= ~a[8];
            a[28] <= ~a[28];
            a[44] <= ~a[44];
            a[22] <= ~a[22];
            #1;
            a[62] <= ~a[62];
            a[9] <= ~a[9];
            a[7] <= ~a[7];
            #1;
            a[18] <= ~a[18];
            #1;
            a[36] <= ~a[36];
            a[1] <= ~a[1];
            a[23] <= ~a[23];
            a[55] <= ~a[55];
            a[59] <= ~a[59];
            a[39] <= ~a[39];
            a[53] <= ~a[53];
            a[6] <= ~a[6];
            a[54] <= ~a[54];
            a[20] <= ~a[20];
            a[27] <= ~a[27];
            #1;
            a[8] <= ~a[8];
            #1;
            a[52] <= ~a[52];
            a[8] <= ~a[8];
            a[36] <= ~a[36];
            a[9] <= ~a[9];
            a[31] <= ~a[31];
            a[20] <= ~a[20];
            #1;
            a[6] <= ~a[6];
            a[45] <= ~a[45];
            a[41] <= ~a[41];
            a[29] <= ~a[29];
            a[13] <= ~a[13];
            #1;
            a[3] <= ~a[3];
            #1;
            a[52] <= ~a[52];
            a[51] <= ~a[51];
            a[61] <= ~a[61];
            a[24] <= ~a[24];
            a[40] <= ~a[40];
            a[55] <= ~a[55];
            a[14] <= ~a[14];
            a[3] <= ~a[3];
            a[18] <= ~a[18];
            a[51] <= ~a[51];
            a[18] <= ~a[18];
            a[20] <= ~a[20];
            a[18] <= ~a[18];
            a[0] <= ~a[0];
            #1;
            a[47] <= ~a[47];
            a[57] <= ~a[57];
            a[32] <= ~a[32];
            a[59] <= ~a[59];
            a[13] <= ~a[13];
            a[0] <= ~a[0];
            a[42] <= ~a[42];
            a[41] <= ~a[41];
            a[59] <= ~a[59];
            a[37] <= ~a[37];
            #1;
            a[56] <= ~a[56];
            a[33] <= ~a[33];
            a[6] <= ~a[6];
            a[18] <= ~a[18];
            a[61] <= ~a[61];
            a[31] <= ~a[31];
            a[29] <= ~a[29];
            a[45] <= ~a[45];
            a[31] <= ~a[31];
            a[12] <= ~a[12];
            a[16] <= ~a[16];
            a[32] <= ~a[32];
            a[7] <= ~a[7];
            a[26] <= ~a[26];
            a[9] <= ~a[9];
            a[32] <= ~a[32];
            a[38] <= ~a[38];
            #1;
            a[61] <= ~a[61];
            a[15] <= ~a[15];
            a[59] <= ~a[59];
            a[58] <= ~a[58];
            a[48] <= ~a[48];
            #1;
            a[54] <= ~a[54];
            a[36] <= ~a[36];
            a[54] <= ~a[54];
            a[63] <= ~a[63];
            a[63] <= ~a[63];
            a[29] <= ~a[29];
            a[59] <= ~a[59];
            #1;
            a[48] <= ~a[48];
            a[38] <= ~a[38];
            a[56] <= ~a[56];
            #1;
            a[15] <= ~a[15];
            #1;
            a[56] <= ~a[56];
            a[43] <= ~a[43];
            #1;
            a[43] <= ~a[43];
            #1;
            a[8] <= ~a[8];
            a[1] <= ~a[1];
            a[25] <= ~a[25];
            a[61] <= ~a[61];
            a[8] <= ~a[8];
            a[50] <= ~a[50];
            a[5] <= ~a[5];
            a[48] <= ~a[48];
            a[14] <= ~a[14];
            a[45] <= ~a[45];
            a[0] <= ~a[0];
            a[55] <= ~a[55];
            a[7] <= ~a[7];
            #1;
            a[0] <= ~a[0];
            a[50] <= ~a[50];
            a[25] <= ~a[25];
            a[53] <= ~a[53];
            #1;
            a[55] <= ~a[55];
            #1;
            a[51] <= ~a[51];
            a[26] <= ~a[26];
            a[31] <= ~a[31];
            a[36] <= ~a[36];
            a[35] <= ~a[35];
            a[16] <= ~a[16];
            a[5] <= ~a[5];
            a[62] <= ~a[62];
            a[40] <= ~a[40];
            a[12] <= ~a[12];
            a[25] <= ~a[25];
            #1;
            a[19] <= ~a[19];
            a[36] <= ~a[36];
            a[21] <= ~a[21];
            a[31] <= ~a[31];
            a[53] <= ~a[53];
            a[1] <= ~a[1];
            #1;
            a[50] <= ~a[50];
            a[22] <= ~a[22];
            a[4] <= ~a[4];
            a[36] <= ~a[36];
            a[12] <= ~a[12];
            #1;
            a[56] <= ~a[56];
            a[3] <= ~a[3];
            a[13] <= ~a[13];
            a[33] <= ~a[33];
            #1;
            a[16] <= ~a[16];
            a[17] <= ~a[17];
            a[1] <= ~a[1];
            #1;
            a[12] <= ~a[12];
            a[52] <= ~a[52];
            #1;
            a[7] <= ~a[7];
            a[3] <= ~a[3];
            #1;
            a[46] <= ~a[46];
            #1;
            a[17] <= ~a[17];
            a[8] <= ~a[8];
            a[49] <= ~a[49];
            a[59] <= ~a[59];
            a[63] <= ~a[63];
            #1;
            a[39] <= ~a[39];
            a[35] <= ~a[35];
            a[6] <= ~a[6];
            a[25] <= ~a[25];
            a[44] <= ~a[44];
            #1;
            a[46] <= ~a[46];
            a[43] <= ~a[43];
            a[12] <= ~a[12];
            a[61] <= ~a[61];
            a[41] <= ~a[41];
            a[54] <= ~a[54];
            a[16] <= ~a[16];
            a[4] <= ~a[4];
            a[57] <= ~a[57];
            a[29] <= ~a[29];
            a[9] <= ~a[9];
            #1;
            a[61] <= ~a[61];
            a[32] <= ~a[32];
            a[37] <= ~a[37];
            a[32] <= ~a[32];
            a[22] <= ~a[22];
            #1;
            a[33] <= ~a[33];
            a[7] <= ~a[7];
            a[6] <= ~a[6];
            #1;
            a[1] <= ~a[1];
            #1;
            a[33] <= ~a[33];
            a[11] <= ~a[11];
            a[17] <= ~a[17];
            #1;
            a[60] <= ~a[60];
            #1;
            a[0] <= ~a[0];
            a[22] <= ~a[22];
            a[3] <= ~a[3];
            a[41] <= ~a[41];
            a[41] <= ~a[41];
            a[8] <= ~a[8];
            a[58] <= ~a[58];
            a[25] <= ~a[25];
            a[22] <= ~a[22];
            #1;
            a[47] <= ~a[47];
            a[1] <= ~a[1];
            a[40] <= ~a[40];
            #1;
            a[48] <= ~a[48];
            a[6] <= ~a[6];
            #1;
            a[26] <= ~a[26];
            a[61] <= ~a[61];
            #1;
            a[54] <= ~a[54];
            a[21] <= ~a[21];
            a[42] <= ~a[42];
            a[12] <= ~a[12];
            a[21] <= ~a[21];
            #1;
            a[33] <= ~a[33];
            a[11] <= ~a[11];
            a[35] <= ~a[35];
            a[26] <= ~a[26];
            a[59] <= ~a[59];
            #1;
            a[16] <= ~a[16];
            a[56] <= ~a[56];
            #1;
            a[33] <= ~a[33];
            #1;
            a[44] <= ~a[44];
            a[60] <= ~a[60];
            a[48] <= ~a[48];
            a[57] <= ~a[57];
            a[28] <= ~a[28];
            a[47] <= ~a[47];
            a[61] <= ~a[61];
            #1;
            a[26] <= ~a[26];
            a[42] <= ~a[42];
            #1;
            a[2] <= ~a[2];
            a[59] <= ~a[59];
            a[8] <= ~a[8];
            #1;
            a[3] <= ~a[3];
            a[21] <= ~a[21];
            a[36] <= ~a[36];
            a[1] <= ~a[1];
            a[41] <= ~a[41];
            a[14] <= ~a[14];
            #1;
            a[50] <= ~a[50];
            a[37] <= ~a[37];
            a[45] <= ~a[45];
            a[7] <= ~a[7];
            a[4] <= ~a[4];
            #1;
            a[25] <= ~a[25];
            a[6] <= ~a[6];
            a[8] <= ~a[8];
            a[53] <= ~a[53];
            a[49] <= ~a[49];
            a[25] <= ~a[25];
            a[18] <= ~a[18];
            a[10] <= ~a[10];
            a[56] <= ~a[56];
            #1;
            a[26] <= ~a[26];
            a[32] <= ~a[32];
            #1;
            a[43] <= ~a[43];
            a[10] <= ~a[10];
            a[21] <= ~a[21];
            a[12] <= ~a[12];
            a[44] <= ~a[44];
            a[16] <= ~a[16];
            #1;
            a[59] <= ~a[59];
            a[12] <= ~a[12];
            #1;
            a[62] <= ~a[62];
            #1;
            a[46] <= ~a[46];
            a[43] <= ~a[43];
            a[26] <= ~a[26];
            a[27] <= ~a[27];
            a[36] <= ~a[36];
            a[62] <= ~a[62];
            a[29] <= ~a[29];
            a[32] <= ~a[32];
            a[46] <= ~a[46];
            a[44] <= ~a[44];
            a[9] <= ~a[9];
            a[3] <= ~a[3];
            a[36] <= ~a[36];
            a[40] <= ~a[40];
            a[61] <= ~a[61];
            a[54] <= ~a[54];
            #1;
            a[20] <= ~a[20];
            a[32] <= ~a[32];
            a[5] <= ~a[5];
            #1;
            a[10] <= ~a[10];
            #1;
            a[23] <= ~a[23];
            a[59] <= ~a[59];
            a[44] <= ~a[44];
            a[20] <= ~a[20];
            #1;
            a[57] <= ~a[57];
            a[34] <= ~a[34];
            a[19] <= ~a[19];
            a[2] <= ~a[2];
            a[31] <= ~a[31];
            a[25] <= ~a[25];
            a[31] <= ~a[31];
            a[31] <= ~a[31];
            #1;
            a[34] <= ~a[34];
            #1;
            a[37] <= ~a[37];
            a[58] <= ~a[58];
            #1;
            a[36] <= ~a[36];
            #1;
            a[29] <= ~a[29];
            a[12] <= ~a[12];
            a[0] <= ~a[0];
            a[18] <= ~a[18];
            a[43] <= ~a[43];
            a[6] <= ~a[6];
            a[24] <= ~a[24];
            a[31] <= ~a[31];
            a[58] <= ~a[58];
            #1;
            a[23] <= ~a[23];
            a[22] <= ~a[22];
            #1;
            a[19] <= ~a[19];
            a[8] <= ~a[8];
            a[56] <= ~a[56];
            #1;
            a[0] <= ~a[0];
            a[51] <= ~a[51];
            a[23] <= ~a[23];
            a[54] <= ~a[54];
            a[38] <= ~a[38];
            #1;
            a[15] <= ~a[15];
            a[61] <= ~a[61];
            #1;
            a[34] <= ~a[34];
            a[50] <= ~a[50];
            a[4] <= ~a[4];
            a[33] <= ~a[33];
            #1;
            a[19] <= ~a[19];
            a[5] <= ~a[5];
            a[19] <= ~a[19];
            a[43] <= ~a[43];
            a[20] <= ~a[20];
            a[40] <= ~a[40];
            a[2] <= ~a[2];
            #1;
            a[38] <= ~a[38];
            a[50] <= ~a[50];
            a[63] <= ~a[63];
            a[60] <= ~a[60];
            #1;
            a[11] <= ~a[11];
            a[5] <= ~a[5];
            a[49] <= ~a[49];
            a[47] <= ~a[47];
            #1;
            a[2] <= ~a[2];
            a[13] <= ~a[13];
            a[41] <= ~a[41];
            #1;
            a[32] <= ~a[32];
            a[61] <= ~a[61];
            a[40] <= ~a[40];
            a[52] <= ~a[52];
            #1;
            a[52] <= ~a[52];
            a[47] <= ~a[47];
            a[31] <= ~a[31];
            a[58] <= ~a[58];
            a[34] <= ~a[34];
            a[43] <= ~a[43];
            a[39] <= ~a[39];
            a[46] <= ~a[46];
            a[61] <= ~a[61];
            a[22] <= ~a[22];
            a[27] <= ~a[27];
            a[0] <= ~a[0];
            a[45] <= ~a[45];
            a[20] <= ~a[20];
            a[47] <= ~a[47];
            a[36] <= ~a[36];
            a[53] <= ~a[53];
            #1;
            a[40] <= ~a[40];
            #1;
            a[29] <= ~a[29];
            #1;
            a[62] <= ~a[62];
            a[53] <= ~a[53];
            #1;
            a[8] <= ~a[8];
            a[1] <= ~a[1];
            a[13] <= ~a[13];
            a[28] <= ~a[28];
            a[50] <= ~a[50];
            a[41] <= ~a[41];
            #1;
            a[48] <= ~a[48];
            a[18] <= ~a[18];
            a[28] <= ~a[28];
            a[13] <= ~a[13];
            a[54] <= ~a[54];
            a[4] <= ~a[4];
            a[2] <= ~a[2];
            a[60] <= ~a[60];
            #1;
            a[17] <= ~a[17];
            a[50] <= ~a[50];
            a[49] <= ~a[49];
            a[52] <= ~a[52];
            a[16] <= ~a[16];
            a[29] <= ~a[29];
            a[19] <= ~a[19];
            a[19] <= ~a[19];
            a[3] <= ~a[3];
            a[32] <= ~a[32];
            a[2] <= ~a[2];
            a[14] <= ~a[14];
            a[12] <= ~a[12];
            a[23] <= ~a[23];
            a[22] <= ~a[22];
            #1;
            a[16] <= ~a[16];
            a[40] <= ~a[40];
            a[50] <= ~a[50];
            a[41] <= ~a[41];
            a[45] <= ~a[45];
            a[19] <= ~a[19];
            a[2] <= ~a[2];
            a[59] <= ~a[59];
            a[0] <= ~a[0];
            a[17] <= ~a[17];
            a[60] <= ~a[60];
            a[54] <= ~a[54];
            a[44] <= ~a[44];
            a[18] <= ~a[18];
            a[13] <= ~a[13];
            a[55] <= ~a[55];
            a[19] <= ~a[19];
            a[0] <= ~a[0];
            a[10] <= ~a[10];
            a[37] <= ~a[37];
            a[19] <= ~a[19];
            #1;
            a[30] <= ~a[30];
            a[29] <= ~a[29];
            a[60] <= ~a[60];
            a[24] <= ~a[24];
            a[9] <= ~a[9];
            a[11] <= ~a[11];
            a[45] <= ~a[45];
            a[59] <= ~a[59];
            a[58] <= ~a[58];
            a[12] <= ~a[12];
            #1;
            a[6] <= ~a[6];
            #1;
            a[59] <= ~a[59];
            a[26] <= ~a[26];
            a[27] <= ~a[27];
            #1;
            a[23] <= ~a[23];
            a[50] <= ~a[50];
            a[30] <= ~a[30];
            a[42] <= ~a[42];
            a[24] <= ~a[24];
            #1;
            a[53] <= ~a[53];
            a[47] <= ~a[47];
            a[47] <= ~a[47];
            a[56] <= ~a[56];
            #1;
            a[19] <= ~a[19];
            #1;
            a[60] <= ~a[60];
            a[32] <= ~a[32];
            a[36] <= ~a[36];
            a[12] <= ~a[12];
            a[1] <= ~a[1];
            a[54] <= ~a[54];
            a[28] <= ~a[28];
            a[54] <= ~a[54];
            #1;
            a[47] <= ~a[47];
            a[3] <= ~a[3];
            a[22] <= ~a[22];
            a[46] <= ~a[46];
            #1;
            a[44] <= ~a[44];
            a[22] <= ~a[22];
            a[26] <= ~a[26];
            a[32] <= ~a[32];
            a[54] <= ~a[54];
            a[6] <= ~a[6];
            a[43] <= ~a[43];
            #1;
            a[40] <= ~a[40];
            a[47] <= ~a[47];
            a[43] <= ~a[43];
            #1;
            a[0] <= ~a[0];
            #1;
            a[25] <= ~a[25];
            a[20] <= ~a[20];
            #1;
            a[8] <= ~a[8];
            a[33] <= ~a[33];
            a[38] <= ~a[38];
            a[25] <= ~a[25];
            #1;
            a[23] <= ~a[23];
            #1;
            a[53] <= ~a[53];
            a[0] <= ~a[0];
            #1;
            a[4] <= ~a[4];
            a[0] <= ~a[0];
            a[7] <= ~a[7];
            a[31] <= ~a[31];
            a[63] <= ~a[63];
            a[45] <= ~a[45];
            a[28] <= ~a[28];
            #1;
            a[43] <= ~a[43];
            #1;
            a[0] <= ~a[0];
            a[39] <= ~a[39];
            #1;
            a[35] <= ~a[35];
            a[47] <= ~a[47];
            a[27] <= ~a[27];
            a[34] <= ~a[34];
            a[48] <= ~a[48];
            a[54] <= ~a[54];
            a[58] <= ~a[58];
            a[15] <= ~a[15];
            #1;
            a[18] <= ~a[18];
            a[48] <= ~a[48];
            a[8] <= ~a[8];
            a[35] <= ~a[35];
            a[14] <= ~a[14];
            a[4] <= ~a[4];
            a[8] <= ~a[8];
            a[17] <= ~a[17];
            a[45] <= ~a[45];
            a[45] <= ~a[45];
            #1;
            a[59] <= ~a[59];
            a[55] <= ~a[55];
            a[61] <= ~a[61];
            a[42] <= ~a[42];
            a[30] <= ~a[30];
            a[54] <= ~a[54];
            #1;
            a[16] <= ~a[16];
            a[23] <= ~a[23];
            #1;
            a[49] <= ~a[49];
            a[11] <= ~a[11];
            a[17] <= ~a[17];
            a[27] <= ~a[27];
            #1;
            a[40] <= ~a[40];
            a[19] <= ~a[19];
            a[18] <= ~a[18];
            a[20] <= ~a[20];
            a[19] <= ~a[19];
            a[1] <= ~a[1];
            a[19] <= ~a[19];
            a[14] <= ~a[14];
            a[62] <= ~a[62];
            a[41] <= ~a[41];
            #1;
            a[53] <= ~a[53];
            #1;
            a[5] <= ~a[5];
            a[58] <= ~a[58];
            a[10] <= ~a[10];
            a[39] <= ~a[39];
            a[59] <= ~a[59];
            a[50] <= ~a[50];
            #1;
            a[29] <= ~a[29];
            a[17] <= ~a[17];
            a[37] <= ~a[37];
            a[42] <= ~a[42];
            a[41] <= ~a[41];
            #1;
            a[6] <= ~a[6];
            a[5] <= ~a[5];
            a[1] <= ~a[1];
            a[59] <= ~a[59];
            #1;
            a[62] <= ~a[62];
            a[36] <= ~a[36];
            #1;
            a[3] <= ~a[3];
            #1;
            a[22] <= ~a[22];
            a[34] <= ~a[34];
            a[34] <= ~a[34];
            a[16] <= ~a[16];
            a[44] <= ~a[44];
            a[57] <= ~a[57];
            #1;
            a[5] <= ~a[5];
            #1;
            a[50] <= ~a[50];
            a[12] <= ~a[12];
            a[25] <= ~a[25];
            a[43] <= ~a[43];
            a[30] <= ~a[30];
            a[1] <= ~a[1];
            #1;
            a[31] <= ~a[31];
            a[11] <= ~a[11];
            a[58] <= ~a[58];
            #1;
            a[0] <= ~a[0];
            a[5] <= ~a[5];
            a[4] <= ~a[4];
            a[49] <= ~a[49];
            #1;
            a[30] <= ~a[30];
            a[27] <= ~a[27];
            a[14] <= ~a[14];
            a[52] <= ~a[52];
            a[55] <= ~a[55];
            a[37] <= ~a[37];
            a[41] <= ~a[41];
            a[10] <= ~a[10];
            a[48] <= ~a[48];
            a[5] <= ~a[5];
            #1;
            a[55] <= ~a[55];
            a[19] <= ~a[19];
            #1;
            a[30] <= ~a[30];
            a[4] <= ~a[4];
            a[45] <= ~a[45];
            a[4] <= ~a[4];
            a[46] <= ~a[46];
            #1;
            a[41] <= ~a[41];
            a[3] <= ~a[3];
            a[22] <= ~a[22];
            #1;
            a[57] <= ~a[57];
            a[5] <= ~a[5];
            a[36] <= ~a[36];
            a[8] <= ~a[8];
            a[45] <= ~a[45];
            a[30] <= ~a[30];
            a[61] <= ~a[61];
            #1;
            a[34] <= ~a[34];
            a[29] <= ~a[29];
            a[22] <= ~a[22];
            a[17] <= ~a[17];
            a[35] <= ~a[35];
            a[30] <= ~a[30];
            a[50] <= ~a[50];
            a[54] <= ~a[54];
            a[17] <= ~a[17];
            a[0] <= ~a[0];
            a[18] <= ~a[18];
            a[59] <= ~a[59];
            a[57] <= ~a[57];
            a[35] <= ~a[35];
            a[9] <= ~a[9];
            a[54] <= ~a[54];
            a[61] <= ~a[61];
            #1;
            a[36] <= ~a[36];
            a[45] <= ~a[45];
            #1;
            a[48] <= ~a[48];
            a[13] <= ~a[13];
            a[58] <= ~a[58];
            #1;
            a[7] <= ~a[7];
            a[23] <= ~a[23];
            a[9] <= ~a[9];
            #1;
            a[12] <= ~a[12];
            a[29] <= ~a[29];
            #1;
            a[29] <= ~a[29];
            a[0] <= ~a[0];
            a[60] <= ~a[60];
            a[0] <= ~a[0];
            a[43] <= ~a[43];
            a[5] <= ~a[5];
            #1;
            a[39] <= ~a[39];
            a[53] <= ~a[53];
            #1;
            a[53] <= ~a[53];
            a[9] <= ~a[9];
            #1;
            a[24] <= ~a[24];
            a[54] <= ~a[54];
            #1;
            a[52] <= ~a[52];
            a[16] <= ~a[16];
            a[45] <= ~a[45];
            a[4] <= ~a[4];
            a[46] <= ~a[46];
            a[55] <= ~a[55];
            #1;
            a[42] <= ~a[42];
            a[43] <= ~a[43];
            #1;
            a[60] <= ~a[60];
            a[52] <= ~a[52];
            a[16] <= ~a[16];
            a[11] <= ~a[11];
            a[36] <= ~a[36];
            a[32] <= ~a[32];
            a[44] <= ~a[44];
            a[59] <= ~a[59];
            #1;
            a[28] <= ~a[28];
            a[4] <= ~a[4];
            a[21] <= ~a[21];
            #1;
            a[3] <= ~a[3];
            #1;
            a[12] <= ~a[12];
            a[44] <= ~a[44];
            a[18] <= ~a[18];
            a[46] <= ~a[46];
            a[63] <= ~a[63];
            a[18] <= ~a[18];
            a[15] <= ~a[15];
            a[42] <= ~a[42];
            a[55] <= ~a[55];
            #1;
            a[59] <= ~a[59];
            a[24] <= ~a[24];
            a[58] <= ~a[58];
            #1;
            a[58] <= ~a[58];
            #1;
            a[37] <= ~a[37];
            a[55] <= ~a[55];
            a[25] <= ~a[25];
            a[20] <= ~a[20];
            #1;
            a[50] <= ~a[50];
            a[6] <= ~a[6];
            a[32] <= ~a[32];
            a[39] <= ~a[39];
            a[46] <= ~a[46];
            a[1] <= ~a[1];
            a[20] <= ~a[20];
            a[30] <= ~a[30];
            a[26] <= ~a[26];
            a[14] <= ~a[14];
            a[50] <= ~a[50];
            a[15] <= ~a[15];
            #1;
            a[59] <= ~a[59];
            a[60] <= ~a[60];
            a[45] <= ~a[45];
            a[18] <= ~a[18];
            #1;
            a[59] <= ~a[59];
            a[29] <= ~a[29];
            #1;
            a[4] <= ~a[4];
            a[22] <= ~a[22];
            #1;
            a[4] <= ~a[4];
            a[5] <= ~a[5];
            a[62] <= ~a[62];
            a[35] <= ~a[35];
            a[46] <= ~a[46];
            #1;
            a[49] <= ~a[49];
            #1;
            a[4] <= ~a[4];
            #1;
            a[42] <= ~a[42];
            a[60] <= ~a[60];
            a[61] <= ~a[61];
            a[11] <= ~a[11];
            a[53] <= ~a[53];
            a[3] <= ~a[3];
            a[32] <= ~a[32];
            a[28] <= ~a[28];
            a[62] <= ~a[62];
            a[31] <= ~a[31];
            a[34] <= ~a[34];
            #1;
            a[33] <= ~a[33];
            #1;
            a[48] <= ~a[48];
            a[13] <= ~a[13];
            a[12] <= ~a[12];
            a[39] <= ~a[39];
            a[54] <= ~a[54];
            a[62] <= ~a[62];
            a[31] <= ~a[31];
            a[29] <= ~a[29];
            a[31] <= ~a[31];
            a[16] <= ~a[16];
            a[17] <= ~a[17];
            a[11] <= ~a[11];
            a[42] <= ~a[42];
            a[43] <= ~a[43];
            a[26] <= ~a[26];
            a[34] <= ~a[34];
            a[61] <= ~a[61];
            a[10] <= ~a[10];
            a[62] <= ~a[62];
            a[44] <= ~a[44];
            a[9] <= ~a[9];
            #1;
            a[36] <= ~a[36];
            a[40] <= ~a[40];
            a[59] <= ~a[59];
            a[6] <= ~a[6];
            a[44] <= ~a[44];
            a[11] <= ~a[11];
            a[12] <= ~a[12];
            a[28] <= ~a[28];
            #1;
            a[4] <= ~a[4];
            a[20] <= ~a[20];
            a[23] <= ~a[23];
            a[28] <= ~a[28];
            a[32] <= ~a[32];
            #1;
            a[5] <= ~a[5];
            #1;
            a[2] <= ~a[2];
            #1;
            a[18] <= ~a[18];
            a[37] <= ~a[37];
            #1;
            a[63] <= ~a[63];
            a[56] <= ~a[56];
            a[42] <= ~a[42];
            a[10] <= ~a[10];
            a[57] <= ~a[57];
            a[56] <= ~a[56];
            #1;
            a[9] <= ~a[9];
            #1;
            a[55] <= ~a[55];
            a[47] <= ~a[47];
            #1;
            a[33] <= ~a[33];
            a[53] <= ~a[53];
            a[12] <= ~a[12];
            a[57] <= ~a[57];
            a[57] <= ~a[57];
            a[58] <= ~a[58];
            a[2] <= ~a[2];
            a[34] <= ~a[34];
            a[8] <= ~a[8];
            a[34] <= ~a[34];
            #1;
            a[27] <= ~a[27];
            a[34] <= ~a[34];
            a[33] <= ~a[33];
            #1;
            a[51] <= ~a[51];
            a[61] <= ~a[61];
            a[42] <= ~a[42];
            #1;
            a[40] <= ~a[40];
            a[21] <= ~a[21];
            a[54] <= ~a[54];
            a[37] <= ~a[37];
            a[9] <= ~a[9];
            a[42] <= ~a[42];
            a[22] <= ~a[22];
            a[1] <= ~a[1];
            a[34] <= ~a[34];
            #1;
            a[56] <= ~a[56];
            a[14] <= ~a[14];
            a[22] <= ~a[22];
            a[61] <= ~a[61];
            a[30] <= ~a[30];
            a[36] <= ~a[36];
            a[57] <= ~a[57];
            a[38] <= ~a[38];
            a[53] <= ~a[53];
            #1;
            a[0] <= ~a[0];
            a[26] <= ~a[26];
            a[30] <= ~a[30];
            a[8] <= ~a[8];
            #1;
            a[27] <= ~a[27];
            a[26] <= ~a[26];
            a[55] <= ~a[55];
            a[28] <= ~a[28];
            a[5] <= ~a[5];
            a[40] <= ~a[40];
            a[40] <= ~a[40];
            a[30] <= ~a[30];
            a[60] <= ~a[60];
            #1;
            a[47] <= ~a[47];
            #1;
            a[27] <= ~a[27];
            a[18] <= ~a[18];
            a[49] <= ~a[49];
            a[16] <= ~a[16];
            #1;
            a[29] <= ~a[29];
            a[22] <= ~a[22];
            a[10] <= ~a[10];
            a[54] <= ~a[54];
            a[46] <= ~a[46];
            #1;
            a[47] <= ~a[47];
            a[46] <= ~a[46];
            a[14] <= ~a[14];
            a[45] <= ~a[45];
            a[10] <= ~a[10];
            a[39] <= ~a[39];
            a[18] <= ~a[18];
            #1;
            a[12] <= ~a[12];
            #1;
            a[59] <= ~a[59];
            a[0] <= ~a[0];
            a[14] <= ~a[14];
            a[60] <= ~a[60];
            #1;
            a[5] <= ~a[5];
            a[40] <= ~a[40];
            a[29] <= ~a[29];
            a[43] <= ~a[43];
            a[26] <= ~a[26];
            a[19] <= ~a[19];
            a[7] <= ~a[7];
            a[53] <= ~a[53];
            a[62] <= ~a[62];
            a[57] <= ~a[57];
            #1;
            a[4] <= ~a[4];
            a[43] <= ~a[43];
            a[51] <= ~a[51];
            a[59] <= ~a[59];
            #1;
            a[30] <= ~a[30];
            a[6] <= ~a[6];
            a[43] <= ~a[43];
            a[53] <= ~a[53];
            a[60] <= ~a[60];
            #1;
            a[32] <= ~a[32];
            #1;
            a[2] <= ~a[2];
            a[21] <= ~a[21];
            #1;
            a[45] <= ~a[45];
            a[46] <= ~a[46];
            a[11] <= ~a[11];
            a[49] <= ~a[49];
            a[27] <= ~a[27];
            a[7] <= ~a[7];
            a[5] <= ~a[5];
            a[15] <= ~a[15];
            a[60] <= ~a[60];
            a[57] <= ~a[57];
            a[53] <= ~a[53];
            #1;
            a[2] <= ~a[2];
            a[56] <= ~a[56];
            #1;
            a[45] <= ~a[45];
            a[8] <= ~a[8];
            a[23] <= ~a[23];
            a[16] <= ~a[16];
            a[32] <= ~a[32];
            a[47] <= ~a[47];
            #1;
            a[5] <= ~a[5];
            #1;
            a[6] <= ~a[6];
            a[47] <= ~a[47];
            a[49] <= ~a[49];
            a[39] <= ~a[39];
            a[36] <= ~a[36];
            a[17] <= ~a[17];
            #1;
            a[47] <= ~a[47];
            #1;
            a[48] <= ~a[48];
            a[45] <= ~a[45];
            a[62] <= ~a[62];
            #1;
            a[37] <= ~a[37];
            #1;
            a[14] <= ~a[14];
            a[52] <= ~a[52];
            a[57] <= ~a[57];
            a[57] <= ~a[57];
            a[7] <= ~a[7];
            a[43] <= ~a[43];
            a[21] <= ~a[21];
            #1;
            a[8] <= ~a[8];
            a[57] <= ~a[57];
            a[18] <= ~a[18];
            #1;
            a[39] <= ~a[39];
            a[14] <= ~a[14];
            #1;
            a[19] <= ~a[19];
            a[45] <= ~a[45];
            a[4] <= ~a[4];
            a[18] <= ~a[18];
            #1;
            a[20] <= ~a[20];
            a[27] <= ~a[27];
            a[9] <= ~a[9];
            a[2] <= ~a[2];
            a[31] <= ~a[31];
            a[8] <= ~a[8];
            a[29] <= ~a[29];
            a[32] <= ~a[32];
            #1;
            a[27] <= ~a[27];
            a[22] <= ~a[22];
            a[1] <= ~a[1];
            a[23] <= ~a[23];
            a[58] <= ~a[58];
            a[24] <= ~a[24];
            a[43] <= ~a[43];
            a[17] <= ~a[17];
            a[14] <= ~a[14];
            #1;
            a[56] <= ~a[56];
            a[47] <= ~a[47];
            a[7] <= ~a[7];
            a[31] <= ~a[31];
            a[19] <= ~a[19];
            a[1] <= ~a[1];
            a[60] <= ~a[60];
            a[12] <= ~a[12];
            a[47] <= ~a[47];
            a[57] <= ~a[57];
            a[63] <= ~a[63];
            a[34] <= ~a[34];
            a[60] <= ~a[60];
            #1;
            a[32] <= ~a[32];
            a[55] <= ~a[55];
            a[27] <= ~a[27];
            a[39] <= ~a[39];
            a[55] <= ~a[55];
            a[22] <= ~a[22];
            a[36] <= ~a[36];
            a[30] <= ~a[30];
            #1;
            a[15] <= ~a[15];
            a[5] <= ~a[5];
            a[12] <= ~a[12];
            a[45] <= ~a[45];
            #1;
            a[13] <= ~a[13];
            a[37] <= ~a[37];
            a[7] <= ~a[7];
            a[18] <= ~a[18];
            a[29] <= ~a[29];
            #1;
            a[32] <= ~a[32];
            a[26] <= ~a[26];
            a[17] <= ~a[17];
            a[54] <= ~a[54];
            a[36] <= ~a[36];
            a[24] <= ~a[24];
            a[49] <= ~a[49];
            a[60] <= ~a[60];
            a[59] <= ~a[59];
            a[27] <= ~a[27];
            a[22] <= ~a[22];
            a[11] <= ~a[11];
            a[17] <= ~a[17];
            #1;
            a[40] <= ~a[40];
            a[57] <= ~a[57];
            a[11] <= ~a[11];
            #1;
            a[35] <= ~a[35];
            a[51] <= ~a[51];
            a[22] <= ~a[22];
            a[2] <= ~a[2];
            a[50] <= ~a[50];
            a[3] <= ~a[3];
            a[53] <= ~a[53];
            a[34] <= ~a[34];
            a[54] <= ~a[54];
            a[15] <= ~a[15];
            a[34] <= ~a[34];
            #1;
            a[41] <= ~a[41];
            #1;
            a[6] <= ~a[6];
            a[31] <= ~a[31];
            a[20] <= ~a[20];
            a[25] <= ~a[25];
            a[45] <= ~a[45];
            a[56] <= ~a[56];
            a[29] <= ~a[29];
            #1;
            a[52] <= ~a[52];
            #1;
            a[29] <= ~a[29];
            a[57] <= ~a[57];
            a[13] <= ~a[13];
            #1;
            a[61] <= ~a[61];
            a[35] <= ~a[35];
            a[18] <= ~a[18];
            a[45] <= ~a[45];
            a[52] <= ~a[52];
            a[20] <= ~a[20];
            #1;
            a[54] <= ~a[54];
            a[43] <= ~a[43];
            a[56] <= ~a[56];
            a[32] <= ~a[32];
            a[14] <= ~a[14];
            a[51] <= ~a[51];
            #1;
            a[10] <= ~a[10];
            a[57] <= ~a[57];
            a[18] <= ~a[18];
            a[62] <= ~a[62];
            #1;
            a[34] <= ~a[34];
            a[11] <= ~a[11];
            #1;
            a[51] <= ~a[51];
            a[63] <= ~a[63];
            #1;
            a[43] <= ~a[43];
            a[7] <= ~a[7];
            a[12] <= ~a[12];
            a[37] <= ~a[37];
            a[6] <= ~a[6];
            a[18] <= ~a[18];
            a[44] <= ~a[44];
            a[11] <= ~a[11];
            a[7] <= ~a[7];
            a[25] <= ~a[25];
            a[8] <= ~a[8];
            a[14] <= ~a[14];
            a[52] <= ~a[52];
            a[24] <= ~a[24];
            a[32] <= ~a[32];
            #1;
            a[21] <= ~a[21];
            a[50] <= ~a[50];
            #1;
            a[21] <= ~a[21];
            a[47] <= ~a[47];
            a[10] <= ~a[10];
            a[26] <= ~a[26];
            a[23] <= ~a[23];
            #1;
            a[26] <= ~a[26];
            a[10] <= ~a[10];
            a[1] <= ~a[1];
            a[39] <= ~a[39];
            #1;
            a[31] <= ~a[31];
            a[40] <= ~a[40];
            a[8] <= ~a[8];
            a[37] <= ~a[37];
            a[49] <= ~a[49];
            a[53] <= ~a[53];
            a[52] <= ~a[52];
            a[30] <= ~a[30];
            a[24] <= ~a[24];
            a[28] <= ~a[28];
            a[9] <= ~a[9];
            a[41] <= ~a[41];
            a[15] <= ~a[15];
            a[60] <= ~a[60];
            #1;
            a[31] <= ~a[31];
            #1;
            a[32] <= ~a[32];
            a[42] <= ~a[42];
            a[60] <= ~a[60];
            a[18] <= ~a[18];
            a[11] <= ~a[11];
            a[37] <= ~a[37];
            #1;
            a[11] <= ~a[11];
            a[25] <= ~a[25];
            a[52] <= ~a[52];
            a[13] <= ~a[13];
            a[62] <= ~a[62];
            a[7] <= ~a[7];
            a[25] <= ~a[25];
            a[17] <= ~a[17];
            #1;
            a[15] <= ~a[15];
            a[10] <= ~a[10];
            a[38] <= ~a[38];
            a[33] <= ~a[33];
            #1;
            a[38] <= ~a[38];
            a[1] <= ~a[1];
            a[60] <= ~a[60];
            #1;
            a[36] <= ~a[36];
            #1;
            a[11] <= ~a[11];
            #1;
            a[47] <= ~a[47];
            a[56] <= ~a[56];
            a[35] <= ~a[35];
            a[42] <= ~a[42];
            a[59] <= ~a[59];
            a[34] <= ~a[34];
            a[43] <= ~a[43];
            a[54] <= ~a[54];
            a[25] <= ~a[25];
            #1;
            a[54] <= ~a[54];
            a[22] <= ~a[22];
            a[14] <= ~a[14];
            a[28] <= ~a[28];
            #1;
            a[22] <= ~a[22];
            a[60] <= ~a[60];
            a[29] <= ~a[29];
            #1;
            a[31] <= ~a[31];
            #1;
            a[57] <= ~a[57];
            a[54] <= ~a[54];
            a[56] <= ~a[56];
            #1;
            a[54] <= ~a[54];
            #1;
            a[2] <= ~a[2];
            a[40] <= ~a[40];
            a[23] <= ~a[23];
            a[30] <= ~a[30];
            a[45] <= ~a[45];
            #1;
            a[51] <= ~a[51];
            a[14] <= ~a[14];
            a[16] <= ~a[16];
            #1;
            a[6] <= ~a[6];
            #1;
            a[28] <= ~a[28];
            a[23] <= ~a[23];
            #1;
            a[33] <= ~a[33];
            a[37] <= ~a[37];
            a[55] <= ~a[55];
            a[56] <= ~a[56];
            a[34] <= ~a[34];
            #1;
            a[49] <= ~a[49];
            a[45] <= ~a[45];
            a[31] <= ~a[31];
            #1;
            a[56] <= ~a[56];
            a[62] <= ~a[62];
            #1;
            a[29] <= ~a[29];
            a[16] <= ~a[16];
            a[11] <= ~a[11];
            a[37] <= ~a[37];
            a[15] <= ~a[15];
            a[47] <= ~a[47];
            a[48] <= ~a[48];
            a[5] <= ~a[5];
            a[42] <= ~a[42];
            #1;
            a[23] <= ~a[23];
            #1;
            a[5] <= ~a[5];
            a[38] <= ~a[38];
            #1;
            a[8] <= ~a[8];
            a[29] <= ~a[29];
            a[8] <= ~a[8];
            a[46] <= ~a[46];
            a[29] <= ~a[29];
            a[60] <= ~a[60];
            a[54] <= ~a[54];
            a[37] <= ~a[37];
            #1;
            a[55] <= ~a[55];
            a[12] <= ~a[12];
            a[5] <= ~a[5];
            a[6] <= ~a[6];
            #1;
            a[2] <= ~a[2];
            #1;
            a[25] <= ~a[25];
            a[7] <= ~a[7];
            a[57] <= ~a[57];
            a[42] <= ~a[42];
            a[13] <= ~a[13];
            a[35] <= ~a[35];
            a[59] <= ~a[59];
            a[53] <= ~a[53];
            a[16] <= ~a[16];
            a[6] <= ~a[6];
            a[50] <= ~a[50];
            a[61] <= ~a[61];
            a[10] <= ~a[10];
            a[19] <= ~a[19];
            a[11] <= ~a[11];
            a[49] <= ~a[49];
            #1;
            a[29] <= ~a[29];
            a[15] <= ~a[15];
            a[14] <= ~a[14];
            a[20] <= ~a[20];
            a[29] <= ~a[29];
            a[47] <= ~a[47];
            a[26] <= ~a[26];
            #1;
            a[48] <= ~a[48];
            a[18] <= ~a[18];
            #1;
            a[46] <= ~a[46];
            a[45] <= ~a[45];
            a[15] <= ~a[15];
            a[21] <= ~a[21];
            #1;
            a[61] <= ~a[61];
            #1;
            a[20] <= ~a[20];
            a[12] <= ~a[12];
            a[0] <= ~a[0];
            a[21] <= ~a[21];
            a[31] <= ~a[31];
            a[42] <= ~a[42];
            a[41] <= ~a[41];
            a[56] <= ~a[56];
            a[17] <= ~a[17];
            a[34] <= ~a[34];
            a[37] <= ~a[37];
            a[34] <= ~a[34];
            a[16] <= ~a[16];
            #1;
            a[11] <= ~a[11];
            a[3] <= ~a[3];
            a[33] <= ~a[33];
            a[34] <= ~a[34];
            #1;
            a[41] <= ~a[41];
            a[54] <= ~a[54];
            a[23] <= ~a[23];
            a[12] <= ~a[12];
            a[3] <= ~a[3];
            a[56] <= ~a[56];
            a[49] <= ~a[49];
            a[47] <= ~a[47];
            #1;
            a[46] <= ~a[46];
            a[62] <= ~a[62];
            a[62] <= ~a[62];
            a[53] <= ~a[53];
            a[55] <= ~a[55];
            a[62] <= ~a[62];
            a[12] <= ~a[12];
            a[55] <= ~a[55];
            a[14] <= ~a[14];
            a[20] <= ~a[20];
            a[4] <= ~a[4];
            a[22] <= ~a[22];
            a[15] <= ~a[15];
            a[29] <= ~a[29];
            a[46] <= ~a[46];
            a[33] <= ~a[33];
            #1;
            a[41] <= ~a[41];
            a[59] <= ~a[59];
            a[57] <= ~a[57];
            a[3] <= ~a[3];
            a[45] <= ~a[45];
            #1;
            a[46] <= ~a[46];
            a[11] <= ~a[11];
            a[26] <= ~a[26];
            a[28] <= ~a[28];
            a[10] <= ~a[10];
            a[63] <= ~a[63];
            #1;
            a[18] <= ~a[18];
            #1;
            a[10] <= ~a[10];
            #1;
            a[45] <= ~a[45];
            a[9] <= ~a[9];
            a[28] <= ~a[28];
            a[14] <= ~a[14];
            a[20] <= ~a[20];
            a[10] <= ~a[10];
            #1;
            a[59] <= ~a[59];
            a[11] <= ~a[11];
            a[52] <= ~a[52];
            #1;
            a[38] <= ~a[38];
            a[39] <= ~a[39];
            #1;
            a[10] <= ~a[10];
            a[10] <= ~a[10];
            a[32] <= ~a[32];
            a[12] <= ~a[12];
            a[1] <= ~a[1];
            a[16] <= ~a[16];
            a[5] <= ~a[5];
            #1;
            a[48] <= ~a[48];
            a[16] <= ~a[16];
            #1;
            a[55] <= ~a[55];
            a[11] <= ~a[11];
            a[46] <= ~a[46];
            a[28] <= ~a[28];
            a[35] <= ~a[35];
            a[48] <= ~a[48];
            a[47] <= ~a[47];
            a[33] <= ~a[33];
            a[39] <= ~a[39];
            a[15] <= ~a[15];
            a[38] <= ~a[38];
            a[24] <= ~a[24];
            a[34] <= ~a[34];
            #1;
            a[16] <= ~a[16];
            a[44] <= ~a[44];
            a[58] <= ~a[58];
            a[56] <= ~a[56];
            a[11] <= ~a[11];
            a[19] <= ~a[19];
            a[8] <= ~a[8];
            #1;
            a[13] <= ~a[13];
            a[14] <= ~a[14];
            a[34] <= ~a[34];
            a[0] <= ~a[0];
            a[22] <= ~a[22];
            a[22] <= ~a[22];
            a[32] <= ~a[32];
            #1;
            a[50] <= ~a[50];
            a[59] <= ~a[59];
            a[14] <= ~a[14];
            a[36] <= ~a[36];
            a[49] <= ~a[49];
            a[43] <= ~a[43];
            a[50] <= ~a[50];
            a[9] <= ~a[9];
            a[54] <= ~a[54];
            a[13] <= ~a[13];
            #1;
            a[5] <= ~a[5];
            a[3] <= ~a[3];
            a[30] <= ~a[30];
            a[51] <= ~a[51];
            a[16] <= ~a[16];
            #1;
            a[32] <= ~a[32];
            a[22] <= ~a[22];
            a[59] <= ~a[59];
            #1;
            a[1] <= ~a[1];
            #1;
            a[13] <= ~a[13];
            #1;
            a[55] <= ~a[55];
            #1;
            a[24] <= ~a[24];
            a[2] <= ~a[2];
            #1;
            a[47] <= ~a[47];
            a[60] <= ~a[60];
            #1;
            a[37] <= ~a[37];
            a[6] <= ~a[6];
            a[48] <= ~a[48];
            a[39] <= ~a[39];
            a[35] <= ~a[35];
            #1;
            a[18] <= ~a[18];
            a[36] <= ~a[36];
            #1;
            a[47] <= ~a[47];
            a[6] <= ~a[6];
            a[54] <= ~a[54];
            a[4] <= ~a[4];
            a[33] <= ~a[33];
            #1;
            a[19] <= ~a[19];
            a[44] <= ~a[44];
            a[49] <= ~a[49];
            #1;
            a[57] <= ~a[57];
            a[20] <= ~a[20];
            a[6] <= ~a[6];
            a[43] <= ~a[43];
            a[3] <= ~a[3];
            a[53] <= ~a[53];
            a[48] <= ~a[48];
            a[52] <= ~a[52];
            a[11] <= ~a[11];
            a[63] <= ~a[63];
            a[21] <= ~a[21];
            #1;
            a[28] <= ~a[28];
            a[7] <= ~a[7];
            a[51] <= ~a[51];
            #1;
            a[9] <= ~a[9];
            #1;
            a[44] <= ~a[44];
            a[3] <= ~a[3];
            #1;
            a[8] <= ~a[8];
            #1;
            a[10] <= ~a[10];
            #1;
            a[57] <= ~a[57];
            a[2] <= ~a[2];
            a[38] <= ~a[38];
            #1;
            a[52] <= ~a[52];
            a[56] <= ~a[56];
            a[63] <= ~a[63];
            #1;
            a[54] <= ~a[54];
            a[45] <= ~a[45];
            #1;
            a[26] <= ~a[26];
            a[33] <= ~a[33];
            a[42] <= ~a[42];
            a[38] <= ~a[38];
            #1;
            a[63] <= ~a[63];
            a[2] <= ~a[2];
            a[8] <= ~a[8];
            a[2] <= ~a[2];
            a[9] <= ~a[9];
            a[44] <= ~a[44];
            a[38] <= ~a[38];
            a[60] <= ~a[60];
            a[23] <= ~a[23];
            a[61] <= ~a[61];
            a[18] <= ~a[18];
            a[46] <= ~a[46];
            a[6] <= ~a[6];
            a[39] <= ~a[39];
            #1;
            a[56] <= ~a[56];
            #1;
            a[46] <= ~a[46];
            a[57] <= ~a[57];
            a[20] <= ~a[20];
            a[49] <= ~a[49];
            #1;
            a[30] <= ~a[30];
            a[41] <= ~a[41];
            #1;
            a[60] <= ~a[60];
            a[58] <= ~a[58];
            #1;
            a[9] <= ~a[9];
            a[49] <= ~a[49];
            a[23] <= ~a[23];
            a[48] <= ~a[48];
            #1;
            a[22] <= ~a[22];
            #1;
            a[22] <= ~a[22];
            a[30] <= ~a[30];
            #1;
            a[9] <= ~a[9];
            a[40] <= ~a[40];
            #1;
            a[52] <= ~a[52];
            a[40] <= ~a[40];
            a[48] <= ~a[48];
            #1;
            a[44] <= ~a[44];
            a[63] <= ~a[63];
            a[63] <= ~a[63];
            a[29] <= ~a[29];
            a[42] <= ~a[42];
            a[42] <= ~a[42];
            a[47] <= ~a[47];
            a[62] <= ~a[62];
            #1;
            a[16] <= ~a[16];
            a[59] <= ~a[59];
            #1;
            a[29] <= ~a[29];
            a[40] <= ~a[40];
            a[28] <= ~a[28];
            a[7] <= ~a[7];
            a[30] <= ~a[30];
            a[19] <= ~a[19];
            #1;
            a[48] <= ~a[48];
            a[34] <= ~a[34];
            a[23] <= ~a[23];
            a[10] <= ~a[10];
            a[36] <= ~a[36];
            a[13] <= ~a[13];
            a[24] <= ~a[24];
            a[7] <= ~a[7];
            a[8] <= ~a[8];
            a[7] <= ~a[7];
            a[9] <= ~a[9];
            a[28] <= ~a[28];
            a[3] <= ~a[3];
            a[49] <= ~a[49];
            a[29] <= ~a[29];
            a[18] <= ~a[18];
            a[6] <= ~a[6];
            a[36] <= ~a[36];
            #1;
            a[41] <= ~a[41];
            a[61] <= ~a[61];
            a[47] <= ~a[47];
            a[57] <= ~a[57];
            #1;
            a[37] <= ~a[37];
            a[5] <= ~a[5];
            a[43] <= ~a[43];
            a[45] <= ~a[45];
            a[12] <= ~a[12];
            a[23] <= ~a[23];
            a[30] <= ~a[30];
            a[13] <= ~a[13];
            a[51] <= ~a[51];
            a[50] <= ~a[50];
            #1;
            a[1] <= ~a[1];
            a[4] <= ~a[4];
            a[44] <= ~a[44];
            a[21] <= ~a[21];
            a[54] <= ~a[54];
            a[56] <= ~a[56];
            a[35] <= ~a[35];
            a[25] <= ~a[25];
            a[35] <= ~a[35];
            a[37] <= ~a[37];
            #1;
            a[55] <= ~a[55];
            a[30] <= ~a[30];
            a[27] <= ~a[27];
            a[6] <= ~a[6];
            a[37] <= ~a[37];
            #1;
            a[30] <= ~a[30];
            a[19] <= ~a[19];
            a[21] <= ~a[21];
            a[35] <= ~a[35];
            a[0] <= ~a[0];
            a[38] <= ~a[38];
            a[10] <= ~a[10];
            #1;
            a[4] <= ~a[4];
            #1;
            a[15] <= ~a[15];
            a[55] <= ~a[55];
            a[33] <= ~a[33];
            a[39] <= ~a[39];
            a[49] <= ~a[49];
            a[35] <= ~a[35];
            #1;
            a[24] <= ~a[24];
            a[9] <= ~a[9];
            a[23] <= ~a[23];
            a[40] <= ~a[40];
            a[3] <= ~a[3];
            a[57] <= ~a[57];
            a[55] <= ~a[55];
            a[2] <= ~a[2];
            a[40] <= ~a[40];
            a[56] <= ~a[56];
            a[4] <= ~a[4];
            a[48] <= ~a[48];
            a[41] <= ~a[41];
            a[21] <= ~a[21];
            #1;
            a[50] <= ~a[50];
            a[52] <= ~a[52];
            a[9] <= ~a[9];
            a[25] <= ~a[25];
            a[32] <= ~a[32];
            a[29] <= ~a[29];
            #1;
            a[18] <= ~a[18];
            #1;
            a[9] <= ~a[9];
            a[11] <= ~a[11];
            a[10] <= ~a[10];
            #1;
            a[59] <= ~a[59];
            a[52] <= ~a[52];
            a[29] <= ~a[29];
            a[28] <= ~a[28];
            a[13] <= ~a[13];
            a[39] <= ~a[39];
            #1;
            a[21] <= ~a[21];
            #1;
            a[33] <= ~a[33];
            a[50] <= ~a[50];
            a[4] <= ~a[4];
            a[1] <= ~a[1];
            a[27] <= ~a[27];
            a[3] <= ~a[3];
            a[2] <= ~a[2];
            a[6] <= ~a[6];
            a[30] <= ~a[30];
            a[0] <= ~a[0];
            a[39] <= ~a[39];
            a[32] <= ~a[32];
            a[20] <= ~a[20];
            a[54] <= ~a[54];
            a[43] <= ~a[43];
            a[63] <= ~a[63];
            a[30] <= ~a[30];
            a[2] <= ~a[2];
            #1;
            a[63] <= ~a[63];
            a[1] <= ~a[1];
            a[16] <= ~a[16];
            #1;
            a[39] <= ~a[39];
            a[1] <= ~a[1];
            #1;
            a[19] <= ~a[19];
            a[61] <= ~a[61];
            a[47] <= ~a[47];
            a[30] <= ~a[30];
            a[21] <= ~a[21];
            a[43] <= ~a[43];
            a[13] <= ~a[13];
            #1;
            a[24] <= ~a[24];
            a[61] <= ~a[61];
            #1;
            a[60] <= ~a[60];
            a[16] <= ~a[16];
            #1;
            a[20] <= ~a[20];
            a[57] <= ~a[57];
            a[17] <= ~a[17];
            a[24] <= ~a[24];
            a[61] <= ~a[61];
            a[3] <= ~a[3];
            a[63] <= ~a[63];
            a[6] <= ~a[6];
            a[20] <= ~a[20];
            #1;
            a[19] <= ~a[19];
            #1;
            a[17] <= ~a[17];
            a[14] <= ~a[14];
            a[48] <= ~a[48];
            a[34] <= ~a[34];
            a[35] <= ~a[35];
            a[37] <= ~a[37];
            a[45] <= ~a[45];
            a[30] <= ~a[30];
            a[25] <= ~a[25];
            #1;
            a[44] <= ~a[44];
            a[50] <= ~a[50];
            #1;
            a[20] <= ~a[20];
            #1;
            a[35] <= ~a[35];
            a[19] <= ~a[19];
            a[51] <= ~a[51];
            a[19] <= ~a[19];
            #1;
            a[43] <= ~a[43];
            a[33] <= ~a[33];
            a[51] <= ~a[51];
            a[58] <= ~a[58];
            #1;
            a[4] <= ~a[4];
            #1;
            a[23] <= ~a[23];
            a[35] <= ~a[35];
            #1;
            a[40] <= ~a[40];
            a[47] <= ~a[47];
            a[3] <= ~a[3];
            a[21] <= ~a[21];
            a[22] <= ~a[22];
            a[30] <= ~a[30];
            a[44] <= ~a[44];
            a[3] <= ~a[3];
            #1;
            a[45] <= ~a[45];
            a[25] <= ~a[25];
            a[35] <= ~a[35];
            a[43] <= ~a[43];
            #1;
            a[49] <= ~a[49];
            a[12] <= ~a[12];
            #1;
            a[28] <= ~a[28];
            a[63] <= ~a[63];
            a[41] <= ~a[41];
            a[35] <= ~a[35];
            a[16] <= ~a[16];
            #1;
            a[12] <= ~a[12];
            a[20] <= ~a[20];
            a[4] <= ~a[4];
            a[35] <= ~a[35];
            a[5] <= ~a[5];
            a[24] <= ~a[24];
            a[49] <= ~a[49];
            a[62] <= ~a[62];
            a[10] <= ~a[10];
            a[62] <= ~a[62];
            a[3] <= ~a[3];
            a[46] <= ~a[46];
            a[14] <= ~a[14];
            a[6] <= ~a[6];
            #1;
            a[3] <= ~a[3];
            a[6] <= ~a[6];
            a[53] <= ~a[53];
            #1;
            a[26] <= ~a[26];
            a[37] <= ~a[37];
            a[36] <= ~a[36];
            a[62] <= ~a[62];
            #1;
            a[26] <= ~a[26];
            a[47] <= ~a[47];
            a[38] <= ~a[38];
            a[39] <= ~a[39];
            #1;
            a[14] <= ~a[14];
            a[56] <= ~a[56];
            a[37] <= ~a[37];
            a[27] <= ~a[27];
            a[30] <= ~a[30];
            a[24] <= ~a[24];
            a[54] <= ~a[54];
            a[32] <= ~a[32];
            a[60] <= ~a[60];
            a[10] <= ~a[10];
            a[17] <= ~a[17];
            a[49] <= ~a[49];
            a[59] <= ~a[59];
            a[12] <= ~a[12];
            a[45] <= ~a[45];
            a[3] <= ~a[3];
            a[49] <= ~a[49];
            a[21] <= ~a[21];
            a[34] <= ~a[34];
            a[58] <= ~a[58];
            a[20] <= ~a[20];
            a[26] <= ~a[26];
            a[16] <= ~a[16];
            a[41] <= ~a[41];
            #1;
            a[61] <= ~a[61];
            a[45] <= ~a[45];
            a[8] <= ~a[8];
            a[2] <= ~a[2];
            a[33] <= ~a[33];
            a[27] <= ~a[27];
            #1;
            a[53] <= ~a[53];
            a[54] <= ~a[54];
            a[5] <= ~a[5];
            a[61] <= ~a[61];
            a[55] <= ~a[55];
            #1;
            a[6] <= ~a[6];
            a[7] <= ~a[7];
            a[57] <= ~a[57];
            a[32] <= ~a[32];
            a[1] <= ~a[1];
            #1;
            a[58] <= ~a[58];
            a[6] <= ~a[6];
            #1;
            a[46] <= ~a[46];
            a[22] <= ~a[22];
            a[53] <= ~a[53];
            a[62] <= ~a[62];
            a[62] <= ~a[62];
            a[33] <= ~a[33];
            a[33] <= ~a[33];
            a[23] <= ~a[23];
            a[22] <= ~a[22];
            a[40] <= ~a[40];
            a[41] <= ~a[41];
            a[20] <= ~a[20];
            #1;
            a[40] <= ~a[40];
            a[14] <= ~a[14];
            a[45] <= ~a[45];
            a[21] <= ~a[21];
            a[19] <= ~a[19];
            a[5] <= ~a[5];
            #1;
            a[51] <= ~a[51];
            a[42] <= ~a[42];
            a[19] <= ~a[19];
            a[6] <= ~a[6];
            a[0] <= ~a[0];
            a[31] <= ~a[31];
            a[1] <= ~a[1];
            #1;
            a[12] <= ~a[12];
            a[13] <= ~a[13];
            a[3] <= ~a[3];
            a[48] <= ~a[48];
            a[4] <= ~a[4];
            a[57] <= ~a[57];
            a[9] <= ~a[9];
            #1;
            a[43] <= ~a[43];
            a[33] <= ~a[33];
            a[57] <= ~a[57];
            a[3] <= ~a[3];
            #1;
            a[9] <= ~a[9];
            #1;
            a[36] <= ~a[36];
            #1;
            a[52] <= ~a[52];
            a[35] <= ~a[35];
            #1;
            a[6] <= ~a[6];
            a[41] <= ~a[41];
            a[11] <= ~a[11];
            a[24] <= ~a[24];
            a[58] <= ~a[58];
            a[17] <= ~a[17];
            a[18] <= ~a[18];
            a[27] <= ~a[27];
            a[32] <= ~a[32];
            a[2] <= ~a[2];
            a[10] <= ~a[10];
            a[1] <= ~a[1];
            a[46] <= ~a[46];
            #1;
            a[0] <= ~a[0];
            a[9] <= ~a[9];
            a[15] <= ~a[15];
            a[51] <= ~a[51];
            #1;
            a[50] <= ~a[50];
            a[31] <= ~a[31];
            a[41] <= ~a[41];
            a[46] <= ~a[46];
            a[1] <= ~a[1];
            #1;
            a[38] <= ~a[38];
            a[11] <= ~a[11];
            a[41] <= ~a[41];
            a[37] <= ~a[37];
            a[21] <= ~a[21];
            a[49] <= ~a[49];
            a[60] <= ~a[60];
            #1;
            a[46] <= ~a[46];
            a[58] <= ~a[58];
            a[27] <= ~a[27];
            a[29] <= ~a[29];
            #1;
            a[24] <= ~a[24];
            a[29] <= ~a[29];
            #1;
            a[19] <= ~a[19];
            a[37] <= ~a[37];
            a[58] <= ~a[58];
            a[35] <= ~a[35];
            a[16] <= ~a[16];
            a[10] <= ~a[10];
            a[28] <= ~a[28];
            #1;
            a[28] <= ~a[28];
            a[0] <= ~a[0];
            a[60] <= ~a[60];
            #1;
            a[0] <= ~a[0];
            a[24] <= ~a[24];
            a[6] <= ~a[6];
            a[25] <= ~a[25];
            a[58] <= ~a[58];
            a[34] <= ~a[34];
            a[19] <= ~a[19];
            a[43] <= ~a[43];
            #1;
            a[43] <= ~a[43];
            #1;
            a[6] <= ~a[6];
            #1;
            a[37] <= ~a[37];
            a[20] <= ~a[20];
            a[2] <= ~a[2];
            #1;
            a[50] <= ~a[50];
            a[31] <= ~a[31];
            a[59] <= ~a[59];
            a[2] <= ~a[2];
            a[63] <= ~a[63];
            a[4] <= ~a[4];
            a[18] <= ~a[18];
            a[37] <= ~a[37];
            a[24] <= ~a[24];
            #1;
            a[3] <= ~a[3];
            a[36] <= ~a[36];
            a[17] <= ~a[17];
            a[61] <= ~a[61];
            a[21] <= ~a[21];
            a[12] <= ~a[12];
            a[15] <= ~a[15];
            a[21] <= ~a[21];
            #1;
            a[50] <= ~a[50];
            #1;
            a[31] <= ~a[31];
            a[20] <= ~a[20];
            a[58] <= ~a[58];
            a[36] <= ~a[36];
            a[5] <= ~a[5];
            a[61] <= ~a[61];
            a[56] <= ~a[56];
            a[58] <= ~a[58];
            #1;
            a[41] <= ~a[41];
            a[56] <= ~a[56];
            a[25] <= ~a[25];
            #1;
            a[24] <= ~a[24];
            a[19] <= ~a[19];
            a[34] <= ~a[34];
            #1;
            a[23] <= ~a[23];
            a[28] <= ~a[28];
            a[21] <= ~a[21];
            a[14] <= ~a[14];
            a[58] <= ~a[58];
            a[53] <= ~a[53];
            a[31] <= ~a[31];
            a[57] <= ~a[57];
            a[27] <= ~a[27];
            #1;
            a[21] <= ~a[21];
            a[1] <= ~a[1];
            a[9] <= ~a[9];
            a[18] <= ~a[18];
            a[48] <= ~a[48];
            a[57] <= ~a[57];
            a[51] <= ~a[51];
            a[44] <= ~a[44];
            a[16] <= ~a[16];
            a[32] <= ~a[32];
            a[15] <= ~a[15];
            a[62] <= ~a[62];
            a[36] <= ~a[36];
            a[8] <= ~a[8];
            a[11] <= ~a[11];
            a[17] <= ~a[17];
            a[14] <= ~a[14];
            a[25] <= ~a[25];
            a[25] <= ~a[25];
            a[19] <= ~a[19];
            a[36] <= ~a[36];
            a[9] <= ~a[9];
            a[62] <= ~a[62];
            a[1] <= ~a[1];
            a[0] <= ~a[0];
            a[0] <= ~a[0];
            a[6] <= ~a[6];
            a[4] <= ~a[4];
            a[17] <= ~a[17];
            a[2] <= ~a[2];
            a[26] <= ~a[26];
            #1;
            a[2] <= ~a[2];
            a[20] <= ~a[20];
            a[24] <= ~a[24];
            a[2] <= ~a[2];
            a[39] <= ~a[39];
            a[40] <= ~a[40];
            a[5] <= ~a[5];
            a[10] <= ~a[10];
            #1;
            a[61] <= ~a[61];
            a[21] <= ~a[21];
            a[57] <= ~a[57];
            #1;
            a[48] <= ~a[48];
            a[55] <= ~a[55];
            a[37] <= ~a[37];
            a[1] <= ~a[1];
            a[35] <= ~a[35];
            a[16] <= ~a[16];
            a[39] <= ~a[39];
            a[41] <= ~a[41];
            a[62] <= ~a[62];
            a[33] <= ~a[33];
            #1;
            a[49] <= ~a[49];
            #1;
            a[32] <= ~a[32];
            a[56] <= ~a[56];
            a[10] <= ~a[10];
            a[0] <= ~a[0];
            a[46] <= ~a[46];
            a[16] <= ~a[16];
            a[33] <= ~a[33];
            a[21] <= ~a[21];
            a[16] <= ~a[16];
            a[47] <= ~a[47];
            a[18] <= ~a[18];
            a[43] <= ~a[43];
            a[46] <= ~a[46];
            #1;
            a[19] <= ~a[19];
            a[38] <= ~a[38];
            a[52] <= ~a[52];
            a[26] <= ~a[26];
            #1;
            a[35] <= ~a[35];
            #1;
            a[0] <= ~a[0];
            a[27] <= ~a[27];
            a[40] <= ~a[40];
            a[19] <= ~a[19];
            a[18] <= ~a[18];
            a[55] <= ~a[55];
            #1;
            a[51] <= ~a[51];
            a[54] <= ~a[54];
            a[63] <= ~a[63];
            a[16] <= ~a[16];
            a[31] <= ~a[31];
            #1;
            a[49] <= ~a[49];
            #1;
            a[59] <= ~a[59];
            #1;
            a[8] <= ~a[8];
            a[40] <= ~a[40];
            a[9] <= ~a[9];
            a[35] <= ~a[35];
            a[27] <= ~a[27];
            a[39] <= ~a[39];
            a[60] <= ~a[60];
            a[27] <= ~a[27];
            #1;
            a[49] <= ~a[49];
            #1;
            a[22] <= ~a[22];
            a[11] <= ~a[11];
            a[57] <= ~a[57];
            a[42] <= ~a[42];
            a[21] <= ~a[21];
            a[47] <= ~a[47];
            a[49] <= ~a[49];
            a[0] <= ~a[0];
            a[58] <= ~a[58];
            a[10] <= ~a[10];
            a[1] <= ~a[1];
            a[19] <= ~a[19];
            a[30] <= ~a[30];
            #1;
            a[50] <= ~a[50];
            a[49] <= ~a[49];
            a[4] <= ~a[4];
            #1;
            a[51] <= ~a[51];
            a[63] <= ~a[63];
            a[14] <= ~a[14];
            a[27] <= ~a[27];
            #1;
            a[6] <= ~a[6];
            a[57] <= ~a[57];
            a[15] <= ~a[15];
            a[27] <= ~a[27];
            a[8] <= ~a[8];
            #1;
            a[48] <= ~a[48];
            a[26] <= ~a[26];
            a[18] <= ~a[18];
            #1;
            a[1] <= ~a[1];
            a[20] <= ~a[20];
            a[43] <= ~a[43];
            #1;
            a[53] <= ~a[53];
            a[14] <= ~a[14];
            a[9] <= ~a[9];
            #1;
            a[19] <= ~a[19];
            a[45] <= ~a[45];
            a[32] <= ~a[32];
            a[18] <= ~a[18];
            a[28] <= ~a[28];
            a[56] <= ~a[56];
            #1;
            a[0] <= ~a[0];
            a[10] <= ~a[10];
            a[51] <= ~a[51];
            a[4] <= ~a[4];
            #1;
            a[53] <= ~a[53];
            a[57] <= ~a[57];
            #1;
            a[35] <= ~a[35];
            a[4] <= ~a[4];
            a[32] <= ~a[32];
            a[37] <= ~a[37];
            a[48] <= ~a[48];
            a[6] <= ~a[6];
            a[40] <= ~a[40];
            a[20] <= ~a[20];
            a[49] <= ~a[49];
            a[26] <= ~a[26];
            a[61] <= ~a[61];
            a[8] <= ~a[8];
            a[48] <= ~a[48];
            a[54] <= ~a[54];
            a[27] <= ~a[27];
            a[50] <= ~a[50];
            a[52] <= ~a[52];
            a[16] <= ~a[16];
            #1;
            a[30] <= ~a[30];
            #1;
            a[57] <= ~a[57];
            a[12] <= ~a[12];
            a[5] <= ~a[5];
            a[40] <= ~a[40];
            #1;
            a[62] <= ~a[62];
            #1;
            a[33] <= ~a[33];
            a[45] <= ~a[45];
            a[29] <= ~a[29];
            a[60] <= ~a[60];
            a[18] <= ~a[18];
            a[28] <= ~a[28];
            a[55] <= ~a[55];
            a[46] <= ~a[46];
            a[32] <= ~a[32];
            a[63] <= ~a[63];
            a[46] <= ~a[46];
            a[49] <= ~a[49];
            a[51] <= ~a[51];
            a[54] <= ~a[54];
            #1;
            a[33] <= ~a[33];
            a[62] <= ~a[62];
            a[39] <= ~a[39];
            a[32] <= ~a[32];
            a[34] <= ~a[34];
            a[19] <= ~a[19];
            a[4] <= ~a[4];
            a[60] <= ~a[60];
            a[49] <= ~a[49];
            a[46] <= ~a[46];
            #1;
            a[9] <= ~a[9];
            #1;
            a[24] <= ~a[24];
            a[48] <= ~a[48];
            a[32] <= ~a[32];
            a[7] <= ~a[7];
            #1;
            a[56] <= ~a[56];
            a[30] <= ~a[30];
            a[13] <= ~a[13];
            a[50] <= ~a[50];
            a[0] <= ~a[0];
            a[49] <= ~a[49];
            a[44] <= ~a[44];
            a[12] <= ~a[12];
            a[22] <= ~a[22];
            a[56] <= ~a[56];
            #1;
            a[26] <= ~a[26];
            a[29] <= ~a[29];
            a[33] <= ~a[33];
            a[2] <= ~a[2];
            a[22] <= ~a[22];
            a[61] <= ~a[61];
            a[54] <= ~a[54];
            a[54] <= ~a[54];
            a[5] <= ~a[5];
            a[54] <= ~a[54];
            a[38] <= ~a[38];
            a[23] <= ~a[23];
            a[48] <= ~a[48];
            #1;
            a[7] <= ~a[7];
            a[47] <= ~a[47];
            a[59] <= ~a[59];
            #1;
            a[26] <= ~a[26];
            a[11] <= ~a[11];
            #1;
            a[42] <= ~a[42];
            a[16] <= ~a[16];
            a[1] <= ~a[1];

        end
        $display ("%x %x %x", a, b, c);
        $finish;
    end
endmodule
